`timescale 1s/1ps
module layer5(clk,reset,x,y,done);
input clk,reset;
output done;
input signed [17:0]x[0:1];
output signed [17:0]y[0:19];
localparam signed [17:0]W[0:39] = {
-59292,-27171,
60279,42319,
21794,14006,
1815,45889,
-25346,-7836,
-6098,-5153,
-4133,69962,
45605,13062,
-81918,58340,
71557,10610,
2930,-62156,
-582,12340,
-631,21824,
26196,43047,
-90353,31071,
-9683,42980,
66576,-42296,
33454,25641,
6868,-18680,
59582,22770
};
localparam signed [35:0]b[0:19] = {
-24130,-48195,50129,34711,50462,54944,-11999,32637,60452,10086,-46241,35623,66240,34456,-44209,54243,45059,55347,66980,11840
};
layer #(18, 36, 15, 2, 20) L5(clk,reset,x,W,b,y,done);
endmodule
